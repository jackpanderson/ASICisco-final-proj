module fixed_point_unit #(parameter TOTAL_BITS = 32,
                          parameter int FRACTIONAL_BITS = 24)
                          (input system_clock, // Main system clock, 96MHZ
                          input rst, // ACTIVE HIGH!!
                          )
endmodule